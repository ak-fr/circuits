// This is the karat_mul module with recursion for project 
// Karatsuba_multiplier_HDL
// Copyright (C) 2020 JC-S
// 
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
// 
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
// GNU General Public License for more details.
// 
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA 02110-1301, USA.

//-----------------------------------------------------------------------------
//
//FILE NAME     : karatsuba_tv.v
//AUTHOR        : JC-S
//FUNCTION      : Main mult module w. recursion for project 
//                Karatsuba_multiplier_HDL
//INITIAL DATE  : 2020/06/29
//VERSION       : 1.1
//CHANGE LOG    : 1.0: initial version.
//
//CHANGE LOG    : 1.1: Use wireal and in the recursion
//-----------------------------------------------------------------------------


module top_module ();
   localparam N = 16;
   localparam log2_N = 4;
   // bit index number 0
   reg [N-1:0] a;
   reg [N-1:0] b;
   reg [2*N - 1:0] ab;
   
   initial begin 
      $display("N = %0d, log2(N) = %0d", N, log2_N);
   end
   
   /*
   stage #(.N(N),
           .log2_N(log2_N),
           .stage_number(2))
   M
     (.inputs(a), 
      .outputs(Ma));
     */ 

   // Instantiate expmob1 and call the instance M
    karat_mult_recursion #(.wI(N),
			   .wO(2*N),
			   .nSTAGE(log2_N))
   AB
     (.iX(a), 
      .iY(Ma),
      .oO(ab));
	
   initial begin // 
      a = 'b1100_0000_0000_0000;
      b = 'b1111_0000_0010_1010;
      // delay of 100 time units
      //#100 a = 'b1111_0000_0000_0000;
      //#100 a = 'b0000_0000_0000_0000;
      // Wait sufficiently enough time
      #10  $display("Time: %0t | a = %d | b = %d | a*b = %d",  $time, a, b, ab);
      #100 $stop; // end of simulation after 1000 units of time
   end

   // Whenever a change of a or Ma occur display both values with the time
   initial begin 
      $monitor("Time: %0t | a = %d | b = %d | a*b = %d",  $time, a, b, ab);
   end


endmodule




module karat_mult_recursion #(parameter wI = 1024,   // Length of the operand iX and iY
			      parameter wO = 2 * wI, // Length of the output 
			      parameter nSTAGE = 10 // log2(wI)
			      )
   (// data IOs
    input wire [wI-1:0]  iX,
    input wire [wI-1:0]  iY,
    output wire [wO-1:0] oO,
    // control IOs
    input wire	 clk,
    input wire	 rst_n,
    input wire	 i_enable,
    output wire o_finish
    );

   localparam wI_pt = wI / 2;

   wire	      finish_p, finish_q, finish_ts;

   wire [wI_pt-1:0] X_hi, X_lo;
   wire [wI_pt-1:0] Y_hi, Y_lo;

   assign  {X_hi, X_lo} = iX;
   assign  {Y_hi, Y_lo} = iY;

   wire   [wI_pt*2-1:0]   p;
   wire [wI_pt*2-1:0]	  q;
   wire [wI_pt:0]	  r;
   wire [wI_pt:0]	  s;

   assign  r = X_hi + X_lo;
   assign  s = Y_hi + Y_lo;

   wire   [wI_pt*2:0]     u;
   assign  u = p + q;

   wire   [wI+1:0]        t;
   wire			  r_hi, s_hi;
   wire [wI_pt-1:0]	  r_lo, s_lo;

   assign  {r_hi, r_lo} = r;
   assign  {s_hi, s_lo} = s;

   wire   [wI-1:0]        t_s;

   generate
      begin: p_eq_Xhi_x_Yhi
	 if(nSTAGE == 1)
	   begin: p_direct_mult
              assign  p = X_hi & Y_hi;
              assign  finish_p = i_enable;
	   end
	 else
	   begin: p_karat_mult
              karat_mult_recursion #(.wI         (wI_pt),
				     .nSTAGE     (nSTAGE-1))
              u_karat_mult_recursion_p (.iX         (X_hi),
					.iY         (Y_hi),
					.oO         (p),
					.clk        (clk),
					.rst_n      (rst_n),
					.i_enable   (i_enable),
					.o_finish   (finish_p)
					);
	   end
      end
   endgenerate

   generate
      begin: q_eq_Xlo_x_Ylo
	 if(nSTAGE == 1)
	   begin: q_direct_mult
              assign  q = X_lo & Y_lo;
              assign  finish_q = i_enable;
	   end
	 else
	   begin: q_karat_mult
              karat_mult_recursion #(
				     .wI         (wI_pt),
				     .nSTAGE     (nSTAGE-1)
				     )
              u_karat_mult_recursion_q (
					.iX         (X_lo),
					.iY         (Y_lo),
					.oO         (q),
					.clk        (clk),
					.rst_n      (rst_n),
					.i_enable   (i_enable),
					.o_finish   (finish_q)
					);
	   end
      end
   endgenerate

   generate
      begin: ts_eq_rlo_x_slo
	 if(nSTAGE == 1)
	   begin: ts_direct_mult
              assign  t_s = r_lo & s_lo;
              assign  finish_ts = i_enable;
	   end
	 else
	   begin: ts_karat_mult
              karat_mult_recursion #(
				     .wI         (wI_pt),
				     .nSTAGE     (nSTAGE-1)
				     )
              u_karat_mult_recursion_ts (
					 .iX         (r_lo),
					 .iY         (s_lo),
					 .oO         (t_s),
					 .clk        (clk),
					 .rst_n      (rst_n),
					 .i_enable   (i_enable),
					 .o_finish   (finish_ts)
					 );
	   end
      end
   endgenerate

   assign t = ((r_hi & s_hi) << wI) + ((r_hi * s_lo + s_hi * r_lo) << wI_pt) + t_s;

   assign oO = (p << wI) + ((t - u) << wI_pt) + q;

   /* -----\/----- EXCLUDED -----\/-----
    // Vivado complains about 
    always  @(posedge clk or negedge rst_n)
    if(!rst_n)
    o_finish    <= 1'b0;
    else
    o_finish    <= finish_p && finish_q && finish_ts;

    -----/\----- EXCLUDED -----/\----- */
endmodule
